module zero16
(
  output wire [15:0] zero16
);

  assign zero16 = 16'b0000_0000_0000_0000;

endmodule